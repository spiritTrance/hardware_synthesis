`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/07 10:58:03
// Design Name: 
// Module Name: mips
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mips(
	input wire clk,rst,
	output wire[31:0] pcF,
	input wire[31:0] instrF,
	output wire [3:0] memwriteM,
	output wire[31:0] aluoutM,writedataM,
	input wire[31:0] readdataM 
);

	datapath dp(
		clk,rst,
		//fetch stage
		pcF,
		instrF,
		//mem stage
		memwriteM,
		aluoutM,writedataM,
		readdataM
	);
	
endmodule
